`ifndef AXI_MST_PKG_SV
`define AXI_MST_PKG_SV

package axi_mst_pkg;
  import uvm_pkg :: *;
  
  `include "uvm_macros.svh"
  
  import axi_mst_agt_pkg :: *;

endpackage

`endif
