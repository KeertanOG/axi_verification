`ifndef AXI_SLV_PKG_SV
`define AXI_SLV_PKG_SV

package axi_slv_pkg;
  import uvm_pkg :: *;
  
  `include "uvm_macros.svh"
  
  import axi_slv_agt_pkg :: *;
  `include "axi_slv_agt_config.sv"
  `include "axi_slv_agent.sv"

endpackage

`endif
