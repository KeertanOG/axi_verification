`ifndef AXI_MST_AGT_PKG_SV
`define AXI_MST_AGT_PKG_SV

package axi_mst_agt_pkg;
  import uvm_pkg :: *;
  
  `include "uvm_macros.svh"
  
  `include "axi_mst_defines.sv"
  `include "axi_mst_agt_config.sv"
  `include "axi_mst_seq_item.sv"
  `include "axi_mst_seqs.sv"  
  `include "axi_mst_seqr.sv"
  `include "axi_mst_mon.sv"
  `include "axi_mst_drv.sv"
  `include "axi_mst_agent.sv"

endpackage

`endif
