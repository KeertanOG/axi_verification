`ifndef AXI_SLV_DEFINES_SV
`define AXI_SLV_DEFINES_SV

`define SV_ADDR_WIDTH 32
`define SV_DATA_WIDTH 32

`endif
