`ifndef AXI_MST_DEFINES_SV
`define AXI_MST_DEFINES_SV

//`define MST_ADDR_WIDTH 32
//`define MST_DATA_WIDTH 32

`endif
