`ifndef AXI_SLV_DEFINES_SV
`define AXI_SLV_DEFINES_SV

//`define SV_ADDR_WIDTH 32
//`define SV_DATA_WIDTH 32

  //enum for operation type
  typedef enum bit[1:0] {SREAD, SWRITE, SRD_WR} sopr_en;

`endif
