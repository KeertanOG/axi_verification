`ifndef AXI_PKG_SV
`define AXI_PKG_SV

package axi_pkg;
  import uvm_pkg :: *;
  
  `include "uvm_macros.svh"
  
  import axi_env_pkg::*;
  `include "axi_base_test.sv"
  `include "axi_mst_inf.sv"
  `include "axi_mst_inf.sv"

endpackage

`endif
